module or_gate(A, B, X);
output X;
input A, B;

  assign X = A || B;
endmodule
