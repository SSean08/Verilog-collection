module full_adder_tb(Sum, Cout);
  output Sum, Cout;

  reg A, B, Cin;
  

  FA(A, B, Cin, Sum, Cout);

  initial
  begin
    A = 0; B = 0; Cin = 0; #10;
    $finish;
  end

endmodule